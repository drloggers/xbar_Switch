//Control Logic
import xbar_pkg::*;


module control_logic
  
  
endmodule 