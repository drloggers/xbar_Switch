// Switching Logic

import xbar_pkg::*;

module switching_logic
  
  
endmodule