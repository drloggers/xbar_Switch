
import xbar_pkg::*;

interface xbar_if(input clk,rst);

logic [ports-1:0]serial_in;
logic [ports-1:0]serial_out;

endinterface
